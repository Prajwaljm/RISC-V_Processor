`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   16:16:52 03/26/2021
// Design Name:   Imm_Gen
// Module Name:   C:/Verilog_projects/COA-Assignment-2-5/Imm_Gen_TEST.v
// Project Name:  COA-Assignment-2-5
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Imm_Gen
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module Imm_Gen_TEST;

	// Inputs
	reg [31:0] I;

	// Outputs
	wire [63:0] imm;

	// Instantiate the Unit Under Test (UUT)
	Imm_Gen uut (
		.imm(imm), 
		.I(I)
	);

	initial begin
		// Initialize Inputs
		I = 0;

		// Wait 100 ns for global reset to finish
		#10;
        
		$monitor($time, "		I=%b		imm=%b", I, imm);
		// Add stimulus here
		
		/*//R-Type instruction		
		#5 I=32'b0000000 00000 00000 000 00000 0110011; //AND //X
		#5 I=32'b0100000 00000 00000 000 00000 0110011; //SUB //X
		#5 I=32'b0100000 00000 00000 010 00000 0110011; //SLT //X
		#5 I=32'b0000000 00000 00000 110 00000 0110011; //OR  //X
		#5 I=32'b0000000 00000 00000 111 00000 0110011; //AND //X
																			  
		//I-Type instructions										  
		#5 I=32'b100000000001 00000 000 00000 0010011; //ADDI //100000000001
		#5 I=32'b000100000100 00000 000 00000 0010011; //ADDI //000100000100
		#5 I=32'b100000000001 00000 011 00000 0010011; //LD   //100000000001
		#5 I=32'b000000110001 00000 011 00000 0010011; //LD   //000000110001
		#5 I=32'b110100000100 00000 011 00000 0010011; //LD   //110100000100
																			  
      //S-Type instructions										  
		#5 I=32'b1000000 00000 00000 011 00001 0100011; //SD  //100000000001
		#5 I=32'b0000001 00000 00000 011 10001 0100011; //SD  //000000110001
		#5 I=32'b1101000 00000 00000 011 00100 0100011; //SD  //110100000100
																			  
		//SB-Type instructions										  
		#5 I=32'b1101000 00000 00000 000 00100 1100011; //BEQ //101010000010
		#5 I=32'b0100010 00000 00000 000 00101 1100011; //BEQ //011000100010*/
		
		//R-Type instruction		
		#5 I=32'b00000000000000000000000000110011; //AND
		#5 I=32'b01000000000000000000000000110011; //SUB
		#5 I=32'b01000000000000000010000000110011; //SLT
		#5 I=32'b00000000000000000110000000110011; //OR 
		#5 I=32'b00000000000000000111000000110011; //AND
																			  
		//I-Type instructions										  
		#5 I=32'b10000000000100000000000000010011; //ADDI
		#5 I=32'b00010000010000000000000000010011; //ADDI
		#5 I=32'b10000000000100000011000000010011; //LD  
		#5 I=32'b00000011000100000011000000010011; //LD  
		#5 I=32'b11010000010000000011000000010011; //LD  
																		  
      //S-Type instructions									  
		#5 I=32'b10000000000000000011000010100011; //SD 
		#5 I=32'b00000010000000000011100010100011; //SD 
		#5 I=32'b11010000000000000011001000100011; //SD 
																		  
		//SB-Type instructions										  
		#5 I=32'b11010000000000000000001001100011; //BEQ
		#5 I=32'b01000100000000000000001011100011; //BEQ
		
		#10 $finish;
	end
      
endmodule

